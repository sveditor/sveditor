`define SOME_DEFINE 1'b1
`define TOP top
`define MUX `TOP.mux

