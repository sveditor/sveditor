
class cls2;

endclass
