
module m;
	property p1;
		a until b;
	endproperty
	property p2;
		a s_until b;
	endproperty
	property p3;
		a until_with b;
	endproperty
	property p4;
		a s_until_with b;
	endproperty	
	
endmodule