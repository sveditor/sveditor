
class xxxx;
endclass
