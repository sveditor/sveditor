class class_2;
endclass
