
`ifndef INCLUDED_CLASS1_SVH
`define INCLUDED_CLASS1_SVH

class class1;

	function new();
	
	endfunction
	
	
	function int get_data();
		return 5;
	endfunction
	
endclass

`endif /* INCLUDED_CLASS1_SVH */
