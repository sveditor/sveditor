
class cls1;
	// Declare a variable named 'a'
	`MY_MACRO(int, a)

endclass
