
`include "defines.svh"

package basic_lib_pkg;
	`include "class1.svh"
	`include "class2.svh"
endpackage
