
package arg_file_multi_include;

	`include "class1.svh"
	`include "class2.svh"
	
endpackage