
package leaf_multimatch_include_pkg;
	`include "cls1.svh"
endpackage