
class pkg2_cls1;

endclass
