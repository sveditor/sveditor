
`ifndef INCLUDED_CLASS2_SVH
`define INCLUDED_CLASS2_SVH

`unknown_define

class class2;

	function new();
	
	endfunction
	
	
	function int get_data();
		return 5;
	endfunction
	
endclass

`endif /* INCLUDED_CLASS2_SVH */
