
module b;
endmodule
