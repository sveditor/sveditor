package pkg;
	`include "../cls1.svh"
	`include "../../incdir/cls2.svh"

endpackage
