/****************************************************************************
 * multi_port_shared_cov_env_pkg.sv
 ****************************************************************************/
`ifndef INCLUDED_multi_port_shared_cov_env_pkg_sv
`define INCLUDED_multi_port_shared_cov_env_pkg_sv

/**
 * Package: multi_port_shared_cov_env_pkg
 * 
 * TODO: Add package documentation
 */
`include "uvm_macros.svh"
package multi_port_shared_cov_env_pkg;
	import uvm_pkg::*;
	import simple_pkt_agent_pkg::*;

	`include "multi_port_shared_cov_env.svh"

endpackage

`endif /* INCLUDED_multi_port_shared_cov_env_pkg_sv */
