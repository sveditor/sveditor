
`ifdef ARG_FILE_DEFINE_PROJ

module arg_file_define_proj;

endmodule

`endif
