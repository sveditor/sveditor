
package pkg1;
	`include "pkg1_cls1.svh"
	`include "pkg1_cls2.svh"
endpackage
