
package sub_package;
	
endpackage
