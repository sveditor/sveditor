

package pkgB;
  class cA;
  endclass
  class cB;
  endclass
endpackage