${file_header}
class ${name}_config extends uvm_object;
	`uvm_object_utils(${name}_config)

endclass

${file_footer}

