
// This file expects that 'pkg1' has already defined macros
package pkg2;
	`include "pkg2_cls1.svh"
	`include "pkg2_cls2.svh"
endpackage