class cls1;
  int		A, B, C, D;

endclass
