

`include "string.svh"
