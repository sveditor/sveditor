

package pkgA;
  class cA;
  endclass
  class cB;
  endclass
endpackage