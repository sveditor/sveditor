

`include "string.svh"
`include "process.svh"
`include "queue.svh"