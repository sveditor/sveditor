
`include "macros.svh"

package root_pkg;

`include "cls1.svh"

endpackage
