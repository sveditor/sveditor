
class pkg1_cls2;

endclass

