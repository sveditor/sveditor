
package root_pkg;
	class root_cls;
	endclass

endpackage

`include "sub_pkg.sv"
