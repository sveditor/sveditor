
`define make_task(name) \
    task name(); \
    endtask