
class my_pkg_file2;
endclass
