
package file1_pkg;
  class cls1;
  endclass

endpackage
