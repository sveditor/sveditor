

package pkgC;
	class cL;
	endclass
endpackage