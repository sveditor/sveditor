
package arg_file_env_var_pkg;

	`include "class1.svh"
	`include "class2.svh"
	
endpackage