
`define PKG1_MACRO1 class
`define PKG1_MACRO2 endclass
class pkg2_cls1;

endclass
