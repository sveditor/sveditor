
// Ensures macros propagate from file to file
package pkg2;
	`include "pkg2_cls1.svh"
	`include "pkg2_cls2.svh"
endpackage