
class cls1;

endclass
