
`define ENABLE_CLASS1
interface top_interface;
	`include "class1.svh"
	`include "class2.svh"
	`include "subdir/class3.svh"
endinterface
