
package pkg_rel_path_include;

	`include "../../target_inc_file.svh"
	
endpackage