
package root;
	`include "./dir1/cls1.svh"
	`include "./dir2/cls2.svh"
endpackage
