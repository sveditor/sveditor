

module m (input a, b);
	a1: assert #0 (a == b);
endmodule	
