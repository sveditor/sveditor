
module `M1_NAME;

endmodule
