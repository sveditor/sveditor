
package my_pkg;
	`include "src/my_pkg_file1.svh"
	`include "src/my_pkg_file2.svh"
	`include "src_sub/my_pkg_file3.svh"
endpackage
