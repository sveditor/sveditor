
module m1;
  reg m1_r1, m1_r2, m1_r3;

endmodule
