
`include "ovm_macros.svh"

class ovm_sequence_utils_macro;
	`ovm_sequencer_utils_begin(ovm_sequence_utils_macro) 
	`ovm_sequencer_utils_end
	
	/** 
	 * Comment
	`ovm_object_utils_begin(TYPE_NAME)
	 */
	
endclass