
package package_cache_non_include_pkg;
	class cls1;
	endclass
	
	class cls2;
	endclass
	
	function void function_1;
	endfunction

endpackage
