
`define MACRO1 A
`define MACRO2 B
