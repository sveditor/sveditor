

	class cS;
	endclass

	