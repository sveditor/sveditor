
class class2_root;

endclass