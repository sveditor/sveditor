
class @name@_driver extends uvm_driver #(@name@_seq_item);

	`uvm_component_utils(@name@_driver)
	
	

endclass