
package top_package;
	
endpackage
