
// Note: bit is a SV keyword, but not a vlog keyword
module bit;

endmodule
