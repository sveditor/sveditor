
`include "simple_proj_macros.svh"
package simple_proj_pkg;
  `include "class1.svh"
  `include "class2.svh"
  `include "class3.svh"
endpackage
