
module `M2_NAME;

endmodule
