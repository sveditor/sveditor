
`define VMM_IN_PACKAGE

`include "vmm.sv"

