
class class1_root;

endclass