
module top(
	input				clk, rst_n,
//	input				rst_n,
	output bit[31:0]	data
	);
	
endmodule