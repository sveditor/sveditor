/****************************************************************************
 * @name@_config.svh
 ****************************************************************************/

class @name@_config extends uvm_object;

endclass
