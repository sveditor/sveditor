
class pkg1_cls1;

endclass

