
package global_field_ref_pkg;
`include "global_field_ref.svh"
endpackage
