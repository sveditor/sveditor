
`include "subdir/defines2.svh"

`define make_function(name) \
    function void name (); \
    endfunction
    
`define accessor_func \
    function void accessor(); \
    endfunction

