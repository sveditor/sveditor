
package basic_lib_pkg;
	`include "class1_2.svh"
	`include "class1.svh"
	`include "class2.svh"
	`include "subdir/class3.svh"
endpackage
