

module sub;

endmodule
