
`ifdef TEST_MODE
module top();
	`include "../xx.svh"
	`include "../../xxx.svh"
	`include "../../../xxxx.svh"
	`include "../../../../xxxxx.svh"
	
endmodule
`endif



