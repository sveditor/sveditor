
class my_pkg_file3;
endclass
