
module arg_file_libpath_2;

endmodule