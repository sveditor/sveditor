
`define ENABLE_CLASS1
interface top_interface;
	`include "class1.SVH"
	`include "class2.SVh"
	`include "subdir/class3.svh"
endinterface
