

package pkgB;
  class cA;
  endclass
  class cB;
  endclass
  `include "cL.svh"
endpackage