
module m;
	property p1;
		##[0:5] done #-# always !rst;
	endproperty	
	
endmodule