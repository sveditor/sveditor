
module arg_file_libpath_1;

endmodule