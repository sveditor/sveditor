
`include "system_tasks.svh"

`include "string.svh"
`include "process.svh"
`include "queue.svh"
`include "array.svh"
`include "covergroup.svh"
