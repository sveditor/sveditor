
module m2;
  reg m2_r1, m2_r2, m2_r3;

endmodule
