
// PKG1_MACRO1 should be 'class'
`PKG1_MACRO1 pkg2_cls2;

`PKG1_MACRO2


