

`include "string.svh"
`include "process.svh"