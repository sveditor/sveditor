
package foo;

import ovm_pkg::*;

class xbus_master_sequencer extends ovm_sequencer #(ovm_sequence_item);
    protected int master_id;

           protected bit m_set_sequences_called = 1;       static protected string m_static_sequences[$];    static protected string m_static_remove_sequences[$];    static function bit add_typewide_sequence(string type_name);      m_static_sequences.push_back(type_name);      return 1;    endfunction   static function bit remove_typewide_sequence(string type_name);      m_static_remove_sequences.push_back(type_name);      for (int i = 0; i < m_static_sequences.size(); i++) begin        if (m_static_sequences[i] == type_name)          m_static_sequences.delete(i);      end      return 1;   endfunction   function void ovm_update_sequence_lib();     if(this.m_set_sequences_called) begin        set_sequences_queue(m_static_sequences);        this.m_set_sequences_called = 0;     end     for (int i = 0; i < m_static_remove_sequences.size(); i++) begin        remove_sequence(m_static_remove_sequences[i]);      end    endfunction             typedef ovm_component_registry #(xbus_master_sequencer,"xbus_master_sequencer") type_id;     static function type_id get_type();       return type_id::get();     endfunction          const static string type_name = "xbus_master_sequencer";     virtual function string get_type_name ();       return type_name;     endfunction          static bit m_fields_checked = 0;     function void m_field_automation (ovm_object tmp_data__,                                       int what__,                                       string str__);     begin       xbus_master_sequencer local_data__;             typedef xbus_master_sequencer ___local_type____;       string string_aa_key;                           if(what__ == OVM_CHECK_FIELDS) begin         if(! ___local_type____::m_fields_checked)           ___local_type____::m_fields_checked=1;         else           return;       end       if(ovm_auto_options_object.recorder != null) begin         ovm_auto_options_object.recorder.scope = m_sc.scope;       end                   super.m_field_automation(tmp_data__, what__, str__);       if(tmp_data__ != null)                          if(!$cast(local_data__, tmp_data__)) return;       if(what__ == OVM_CHECK_FIELDS) begin         super.m_delete_field_array();       end 
            begin    if(what__==OVM_CHECK_FIELDS) m_do_field_check("master_id");    m_sc.scope.set_arg("master_id");       begin      int r__;      if((what__ == OVM_PRINT) && (((OVM_ALL_ON)&OVM_NOPRINT) == 0) && (ovm_radix_enum'((OVM_ALL_ON)&OVM_RADIX) == OVM_ENUM) &&          (ovm_auto_options_object.printer.knobs.print_fields == 1)) begin        $swrite(m_sc.stringv, "%0d", master_id);        ovm_auto_options_object.printer.print_generic("master_id", "enum",            $bits(master_id), m_sc.stringv);      end      else if((what__ == OVM_RECORD) && (((OVM_ALL_ON)&OVM_NORECORD) == 0) && (ovm_radix_enum'((OVM_ALL_ON)&OVM_RADIX) == OVM_ENUM))      begin        $swrite(m_sc.stringv, "%0d", master_id);        ovm_auto_options_object.recorder.record_string("master_id",m_sc.stringv);      end      else if(tmp_data__!=null) begin        if($cast(local_data__, tmp_data__)) begin          r__ = m_do_data("master_id", master_id, local_data__.master_id, what__, $bits(master_id), OVM_ALL_ON);        end      end      else begin        if(what__ != OVM_COMPARE && what__ != OVM_COPY) begin          r__ = m_do_data("master_id", master_id, 0, what__, $bits(master_id), OVM_ALL_ON);        end      end      if((what__ == OVM_COMPARE) && r__) begin        if(ovm_radix_enum'((OVM_ALL_ON)&OVM_RADIX) == OVM_ENUM) begin          if(local_data__!=null) begin               begin      ovm_comparer comparer;      comparer = ovm_auto_options_object.comparer;      if(comparer==null) comparer = ovm_default_comparer;      comparer.result++;                     $swrite(comparer.miscompares,"%s%s: lhs = %0d : rhs = %0d\n",         comparer.miscompares, comparer.scope.get_arg(), master_id, local_data__.master_id );    end          end          else begin               begin      ovm_comparer comparer;      comparer = ovm_auto_options_object.comparer;      if(comparer==null) comparer = ovm_default_comparer;      comparer.result++;                     $swrite(comparer.miscompares,"%s%s: lhs = %0d : rhs = %0d\n",         comparer.miscompares, comparer.scope.get_arg(), master_id, 0 );    end          end        end      end    end        if(ovm_object::m_do_set (str__, "master_id", master_id, what__, OVM_ALL_ON)) begin      m_sc.scope.up(null);      return;    end    m_sc.scope.unset_arg("master_id");    end
              end     endfunction

endclass

endpackage


