
// PKG1_MACRO1 should be 'class'
`PKG1_MACRO1 pkg1_cls2;

`PKG1_MACRO2


