
class p2_c;

endclass
