
class my_cls2;

endclass
