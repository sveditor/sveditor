
class class3;
endclass