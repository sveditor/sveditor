

`define make_function(name) \
    function void name(); \
    endfunction

