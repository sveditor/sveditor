
module a;
endmodule
