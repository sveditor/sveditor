
module fsm();
	function bit f (int a, int b);
		// ...
		a1: assert #0 (a == b);
		// ...
	endfunction

	always_comb begin : b1
		some_stuff = f(x,y); // ? ...
		// ...
	end
	
	always_comb begin : b2
		other_stuff = f(z,w); // ? ...
		// ...
	end
endmodule