
package sub_pkg;
	`include "sub_cls.svh"

endpackage
