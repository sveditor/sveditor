
`define ENABLE_CLASS1
module top_module;
	`include "class1.svh"
	`include "class2.svh"
	`include "subdir/class3.svh"
endmodule
