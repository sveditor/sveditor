
class cL;
endclass
