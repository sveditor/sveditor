/****************************************************************************
 * ${name}_tb.sv
 ****************************************************************************/

/**
 * Module: ${name}_tb
 * 
 * TODO: Add module documentation
 */
`include "uvm_macros.svh"
module ${name}_tb;
	import uvm_pkg::*;
	import ${name}_tests_pkg::*;
	
	initial begin
		run_test();
	end

endmodule

