module top;

endmodule
