

class simple_agent_test_seq_item extends simple_seq_item;
	`uvm_object_utils(simple_agent_test_seq_item)
	
	int					A;
	int					B;
	
endclass
