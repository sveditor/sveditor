
`define ovm_object_utils(cls)