
package sub_sub_package;
	
endpackage
