
class cls2;
  int D, E, F, G;
  cls1 c1_A, c1_B, c1_C;
endclass
