/********************************************************************
 * @name@_agent.svh
 *
 ********************************************************************/

class @name@_agent extends uvm_agent;

endclass