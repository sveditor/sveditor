
package leaf_multimatch_include_pkg;
	`include "my_cls1.svh"
endpackage