class xxxxx;
endclass
