
class xx;
	
endclass