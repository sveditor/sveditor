
class my_pkg_file1;
endclass
