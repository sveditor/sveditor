
class class2;

endclass