

	class cR;
	endclass

	