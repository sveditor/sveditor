
class class1;

endclass