
package package_cache_include_pkg;
	`include "cls1.svh"

	`include "cls2.svh"	
	
endpackage
