
`ifndef INCLUDED_CLASS3_SVH
`define INCLUDED_CLASS3_SVH

class class3;

	function new();
	
	endfunction
	
	
	function int get_data();
		return 5;
	endfunction
	
endclass

`endif /* INCLUDED_CLASS3_SVH */
