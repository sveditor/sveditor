
class cls_top;
  cls2 c2_A, c2_B, c2_C;
endclass
