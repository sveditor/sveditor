
package pkg;
	`include "cls1.svh"
	`include "cls2.svh"
	`include "cls_top.svh"
endpackage
