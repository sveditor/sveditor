

package src_collection_data_pkg;
	`include "cls1.svh"
	`include "cls2.svh"
endpackage
