
class xxx;
endclass