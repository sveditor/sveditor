
class class2_dir2;

endclass