
class p1_c;

endclass
