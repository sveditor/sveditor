class class_1;
endclass
