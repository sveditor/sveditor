
module m;
	property p2;
		##[0:5] done #=# always !rst;
	endproperty	
	
endmodule
