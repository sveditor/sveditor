
module expected_module;

endmodule

`ifndef EXCLUDE_DEFINED
module arg_file_define_proj;

endmodule
`endif /* EXCLUDE_DEFINED */

