
`define MY_MACRO(t,n) \
  t			n;