/****************************************************************************
 * target_inc_file.svh
 *
 * 
 ****************************************************************************/

class target_inc;
	int m_data;
endclass
