
class global_field_cls;
	int		AA;
	int		AB;
	int		BB;
	int		BA;
endclass

const global_field_cls field_cls = global_field_cls::get();

