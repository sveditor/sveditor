
class class1_dir1;

endclass