
class my_cls1;

endclass
