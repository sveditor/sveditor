
class sub_cls;
endclass
