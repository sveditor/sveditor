
`define M1_NAME m1
`define M2_NAME m2

module top;

	m1		m1_i();
	m2		m2_i();

endmodule
