
`ifndef INCLUDED_CLASS1_SVH    
`define INCLUDED_CLASS1_SVH

class class1;

typedef struct {
int a;
int b;
} foobar;

	/****************************************************************
	 * new()
	 ****************************************************************/
virtual	function new(int a, 
		int b);
	
foo = boolean'(get_bit());
	endfunction
	
	
	function int get_data();
			/**********************************
			 			*
		*
		**********************************/
		if (foobar) begin
			foo = 2;
				if (foo2) begin
						foo2 = 2;
					end // end1
		end // end2
		
		if (foobar)
		foo3 = 3;
		
	while (true) begin
	foobar = 5;
	end
	
	
	
		return 'h5;
	endfunction
	
	
endclass

`endif /* INCLUDED_CLASS1_SVH */
