
`define ENABLE_CLASS1
program top_program;
	`include "class1.svh"
	`include "class2.svh"
	`include "subdir/class3.svh"
endprogram
