
class class1_dir2;

endclass